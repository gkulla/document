library IEEE;
USE IEEE.std_logic_1164.all;


ENTITY Multiplier IS
port ( A, B, C, D: in std_logic;
   out0,out1,out2,out3: out std_logic
      );
END Multiplier;

Architecture Struct OF Multiplier IS
Begin
--F0 = A B C D;
--F1 = A B' C  + A C D';
--F2 = A' B C  + A B' D + A C' D + B C D';
--F3 = B D;
out0 <= A and B and C and D;
out1 <= (A and not B and C)or(A and C and not D);
out2 <= (not A and B and C)or(A and not B and D)or(A and not C and D)or(B and C and not D);
out3 <= B and D;
END Struct;