library IEEE;
use IEEE.std_logic_1164.all;

ENTITY decoder_tre_to_eight IS
port ( a : in std_logic_vector(1 downto 0);
       en: in std_logic;
       f : out std_logic_vector(7 downto 0)
      );
END decoder_tre_to_eight;

Architecture Behav OF decoder_tre_to_eight IS
BEGIN
	Process(en, a)
	Begin
	f <= "00000000"; 
		if(en = '0') then
				 case a is
				 when "00" => f(0) <= '1';--not a(1) and not a(0);
				 when "01" => f(1) <= '1';--not a(1) and  a(0);
				 when "10" => f(2) <= '1';--    a(1) and not a(0);
				 when "11" => f(3) <= '1';--    a(1) and  a(0);
				 when others => f <= "00000000";
				 end case;
		 else
				 case a is 
				 when "00" => f(4) <= '1';--not a(1) and not a(0);
				 when "01" => f(5) <= '1';--not a(1) and  a(0);
				 when "10" => f(6) <= '1';--    a(1) and not a(0);
				 when "11" => f(7) <= '1';--    a(1) and  a(0);
				 when others => f <= "00000000";
			END case;
		END IF;
	END PROCESS;
END Behav;